--
--
--lol im not commenting the og code 
--
--
--
--
LIBRARY ieee;

USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;


ENTITY skip IS
    PORT (
        rng_lo_input : IN UNSIGNED(63 DOWNTO 0);
        rng_hi_input : IN UNSIGNED(63 DOWNTO 0);
        rng_lo_output : OUT UNSIGNED(63 DOWNTO 0);
        rng_hi_output : OUT UNSIGNED(63 DOWNTO 0)
    );
END skip;
ARCHITECTURE arch OF skip IS
    BEGIN

rng_lo_output(0) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(6) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(22) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(49) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(11) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(38) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(1) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(13) XOR rng_lo_input(15) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(22) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(35) XOR rng_lo_input(38) XOR rng_lo_input(41) XOR rng_lo_input(44) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(60) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(47) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(56) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(63);
rng_lo_output(2) <= rng_lo_input(0) XOR rng_lo_input(2) XOR rng_lo_input(6) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(37) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(14) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(21) XOR rng_hi_input(23) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(30) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(53) XOR rng_hi_input(59) XOR rng_hi_input(63);
rng_lo_output(3) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(7) XOR rng_lo_input(9) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(43) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(63) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(7) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(17) XOR rng_hi_input(20) XOR rng_hi_input(23) XOR rng_hi_input(25) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(36) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(56) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(4) <= rng_lo_input(1) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(39) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(54) XOR rng_lo_input(57) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(6) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(15) XOR rng_hi_input(20) XOR rng_hi_input(23) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(39) XOR rng_hi_input(42) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(61);
rng_lo_output(5) <= rng_lo_input(1) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(29) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(37) XOR rng_lo_input(45) XOR rng_lo_input(50) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(4) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(15) XOR rng_hi_input(19) XOR rng_hi_input(23) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(48) XOR rng_hi_input(51) XOR rng_hi_input(55) XOR rng_hi_input(57) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(6) <= rng_lo_input(1) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(8) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(11) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(38) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(63);
rng_lo_output(7) <= rng_lo_input(0) XOR rng_lo_input(5) XOR rng_lo_input(8) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(40) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(58) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(4) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(47) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(62);
rng_lo_output(8) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(9) XOR rng_lo_input(12) XOR rng_lo_input(17) XOR rng_lo_input(21) XOR rng_lo_input(25) XOR rng_lo_input(27) XOR rng_lo_input(29) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(56) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_hi_input(0) XOR rng_hi_input(2) XOR rng_hi_input(6) XOR rng_hi_input(12) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(19) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(30) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(42) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(59);
rng_lo_output(9) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(14) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(60) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(4) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(15) XOR rng_hi_input(19) XOR rng_hi_input(24) XOR rng_hi_input(27) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(46) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(53) XOR rng_hi_input(55) XOR rng_hi_input(59);
rng_lo_output(10) <= rng_lo_input(0) XOR rng_lo_input(2) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(2) XOR rng_hi_input(4) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(11) <= rng_lo_input(0) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(20) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(27) XOR rng_lo_input(29) XOR rng_lo_input(31) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(43) XOR rng_lo_input(45) XOR rng_lo_input(55) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(5) XOR rng_hi_input(9) XOR rng_hi_input(13) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(22) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(43) XOR rng_hi_input(47) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(56) XOR rng_hi_input(59) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(12) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(31) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(45) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(21) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(13) <= rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(15) XOR rng_lo_input(19) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(26) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(41) XOR rng_lo_input(48) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(62) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(12) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(53) XOR rng_hi_input(55) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(14) <= rng_lo_input(0) XOR rng_lo_input(2) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(48) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(62) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(10) XOR rng_hi_input(13) XOR rng_hi_input(21) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(30) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(38) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(61);
rng_lo_output(15) <= rng_lo_input(0) XOR rng_lo_input(4) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(15) XOR rng_lo_input(17) XOR rng_lo_input(21) XOR rng_lo_input(24) XOR rng_lo_input(37) XOR rng_lo_input(40) XOR rng_lo_input(44) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(40) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(56) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(16) <= rng_lo_input(2) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(42) XOR rng_lo_input(45) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(2) XOR rng_hi_input(4) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(12) XOR rng_hi_input(14) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(28) XOR rng_hi_input(30) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(37) XOR rng_hi_input(42) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(60) XOR rng_hi_input(63);
rng_lo_output(17) <= rng_lo_input(0) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(58) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(7) XOR rng_hi_input(10) XOR rng_hi_input(16) XOR rng_hi_input(19) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(30) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(38) XOR rng_hi_input(41) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(56) XOR rng_hi_input(61) XOR rng_hi_input(63);
rng_lo_output(18) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(7) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(17) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(29) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(43) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(62) XOR rng_hi_input(0) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(11) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(35) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(53) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(60) XOR rng_hi_input(62);
rng_lo_output(19) <= rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(12) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(25) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(43) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(63) XOR rng_hi_input(1) XOR rng_hi_input(6) XOR rng_hi_input(10) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(35) XOR rng_hi_input(38) XOR rng_hi_input(41) XOR rng_hi_input(43) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60);
rng_lo_output(20) <= rng_lo_input(0) XOR rng_lo_input(3) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(40) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(1) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(31) XOR rng_hi_input(36) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(58) XOR rng_hi_input(62);
rng_lo_output(21) <= rng_lo_input(1) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(15) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(48) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(60) XOR rng_hi_input(0) XOR rng_hi_input(3) XOR rng_hi_input(8) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(13) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(36) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(49) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(63);
rng_lo_output(22) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(22) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(37) XOR rng_lo_input(40) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(6) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(16) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(30) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(55) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(23) <= rng_lo_input(1) XOR rng_lo_input(9) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(23) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(35) XOR rng_hi_input(38) XOR rng_hi_input(43) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(59);
rng_lo_output(24) <= rng_lo_input(0) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(18) XOR rng_lo_input(21) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(39) XOR rng_lo_input(44) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(10) XOR rng_hi_input(13) XOR rng_hi_input(15) XOR rng_hi_input(21) XOR rng_hi_input(23) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(35) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(47) XOR rng_hi_input(50) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_lo_output(25) <= rng_lo_input(1) XOR rng_lo_input(3) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(47) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(54) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(30) XOR rng_hi_input(34) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(45) XOR rng_hi_input(47) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(57) XOR rng_hi_input(61) XOR rng_hi_input(63);
rng_lo_output(26) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(22) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(41) XOR rng_lo_input(44) XOR rng_lo_input(50) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(8) XOR rng_hi_input(12) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(59) XOR rng_hi_input(61);
rng_lo_output(27) <= rng_lo_input(0) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(13) XOR rng_hi_input(15) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(30) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(56) XOR rng_hi_input(60) XOR rng_hi_input(63);
rng_lo_output(28) <= rng_lo_input(2) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(27) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(36) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(7) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(25) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(46) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(62);
rng_lo_output(29) <= rng_lo_input(1) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(26) XOR rng_lo_input(29) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(41) XOR rng_lo_input(43) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(11) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(23) XOR rng_hi_input(25) XOR rng_hi_input(28) XOR rng_hi_input(30) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(44) XOR rng_hi_input(49) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_lo_output(30) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(13) XOR rng_lo_input(15) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(39) XOR rng_lo_input(41) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(58) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(6) XOR rng_hi_input(10) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(55) XOR rng_hi_input(58) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(31) <= rng_lo_input(1) XOR rng_lo_input(4) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(46) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(12) XOR rng_hi_input(14) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(55) XOR rng_hi_input(57) XOR rng_hi_input(60) XOR rng_hi_input(61);
rng_lo_output(32) <= rng_lo_input(0) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(15) XOR rng_lo_input(17) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(23) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(56) XOR rng_hi_input(59) XOR rng_hi_input(61) XOR rng_hi_input(63);
rng_lo_output(33) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(15) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(44) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(23) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(37) XOR rng_hi_input(41) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(58) XOR rng_hi_input(61);
rng_lo_output(34) <= rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(41) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(49) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_hi_input(0) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(15) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(38) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(62);
rng_lo_output(35) <= rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(13) XOR rng_lo_input(15) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(29) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(53) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(23) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(56) XOR rng_hi_input(58) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(36) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(41) XOR rng_lo_input(43) XOR rng_lo_input(45) XOR rng_lo_input(48) XOR rng_lo_input(51) XOR rng_lo_input(54) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(60) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(12) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(26) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(38) XOR rng_hi_input(42) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60);
rng_lo_output(37) <= rng_lo_input(0) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(17) XOR rng_lo_input(20) XOR rng_lo_input(24) XOR rng_lo_input(28) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(54) XOR rng_lo_input(59) XOR rng_lo_input(62) XOR rng_hi_input(0) XOR rng_hi_input(4) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(15) XOR rng_hi_input(20) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(47) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(61) XOR rng_hi_input(63);
rng_lo_output(38) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(10) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(21) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(31) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(46) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(19) XOR rng_hi_input(23) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(44) XOR rng_hi_input(46) XOR rng_hi_input(48) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_lo_output(39) <= rng_lo_input(0) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(38) XOR rng_lo_input(40) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(3) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(11) XOR rng_hi_input(13) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(38) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(55) XOR rng_hi_input(59) XOR rng_hi_input(63);
rng_lo_output(40) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(10) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(41) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(21) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(32) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(47) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(63);
rng_lo_output(41) <= rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(11) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(49) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(60) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(17) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(47) XOR rng_hi_input(53) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(57);
rng_lo_output(42) <= rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(19) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(45) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(28) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(44) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_lo_output(43) <= rng_lo_input(2) XOR rng_lo_input(5) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(15) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(46) XOR rng_lo_input(52) XOR rng_lo_input(55) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(54) XOR rng_hi_input(58) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(63);
rng_lo_output(44) <= rng_lo_input(0) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(36) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(43) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(51) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(30) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(45) <= rng_lo_input(0) XOR rng_lo_input(2) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(37) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(11) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(21) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(30) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(56) XOR rng_hi_input(60) XOR rng_hi_input(63);
rng_lo_output(46) <= rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(31) XOR rng_lo_input(34) XOR rng_lo_input(37) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(56) XOR rng_lo_input(60) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(28) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(62);
rng_lo_output(47) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(49) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(58) XOR rng_hi_input(0) XOR rng_hi_input(2) XOR rng_hi_input(4) XOR rng_hi_input(7) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(30) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(45) XOR rng_hi_input(48) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_lo_output(48) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(15) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(49) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_hi_input(0) XOR rng_hi_input(2) XOR rng_hi_input(4) XOR rng_hi_input(7) XOR rng_hi_input(11) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(23) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(47) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(60) XOR rng_hi_input(63);
rng_lo_output(49) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(25) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(39) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(58) XOR rng_lo_input(60) XOR rng_hi_input(0) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(33) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(44) XOR rng_hi_input(47) XOR rng_hi_input(50) XOR rng_hi_input(53) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(58) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(63);
rng_lo_output(50) <= rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(7) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(27) XOR rng_lo_input(29) XOR rng_lo_input(35) XOR rng_lo_input(38) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(56) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(0) XOR rng_hi_input(4) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(29) XOR rng_hi_input(34) XOR rng_hi_input(37) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(59);
rng_lo_output(51) <= rng_lo_input(0) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(10) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(27) XOR rng_lo_input(29) XOR rng_lo_input(31) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(43) XOR rng_lo_input(50) XOR rng_lo_input(53) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(60) XOR rng_lo_input(63) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(10) XOR rng_hi_input(13) XOR rng_hi_input(15) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(38) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(53) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(52) <= rng_lo_input(2) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(41) XOR rng_lo_input(45) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(57) XOR rng_lo_input(60) XOR rng_lo_input(63) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(17) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(32) XOR rng_hi_input(37) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(49) XOR rng_hi_input(53) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_lo_output(53) <= rng_lo_input(0) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(21) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(39) XOR rng_lo_input(41) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(56) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(13) XOR rng_hi_input(16) XOR rng_hi_input(19) XOR rng_hi_input(23) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(30) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(48) XOR rng_hi_input(50) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(63);
rng_lo_output(54) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(9) XOR rng_lo_input(11) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(49) XOR rng_lo_input(52) XOR rng_lo_input(58) XOR rng_lo_input(60) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(22) XOR rng_hi_input(25) XOR rng_hi_input(30) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(45) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(62);
rng_lo_output(55) <= rng_lo_input(2) XOR rng_lo_input(4) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(13) XOR rng_lo_input(15) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(22) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(42) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(59) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(53) XOR rng_hi_input(55) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(61);
rng_lo_output(56) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(15) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(28) XOR rng_lo_input(32) XOR rng_lo_input(37) XOR rng_lo_input(40) XOR rng_lo_input(46) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(58) XOR rng_lo_input(61) XOR rng_hi_input(0) XOR rng_hi_input(2) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(23) XOR rng_hi_input(29) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(43) XOR rng_hi_input(47) XOR rng_hi_input(51) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_lo_output(57) <= rng_lo_input(0) XOR rng_lo_input(4) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(38) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(46) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(2) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(53) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(63);
rng_lo_output(58) <= rng_lo_input(0) XOR rng_lo_input(2) XOR rng_lo_input(4) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(11) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(20) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(35) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(40) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(21) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(36) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(50) XOR rng_hi_input(53) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60);
rng_lo_output(59) <= rng_lo_input(1) XOR rng_lo_input(3) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(26) XOR rng_lo_input(29) XOR rng_lo_input(33) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(61) XOR rng_hi_input(0) XOR rng_hi_input(4) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(10) XOR rng_hi_input(13) XOR rng_hi_input(15) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(44) XOR rng_hi_input(46) XOR rng_hi_input(49) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(60) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(60) <= rng_lo_input(0) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(34) XOR rng_lo_input(37) XOR rng_lo_input(40) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(60) XOR rng_hi_input(0) XOR rng_hi_input(3) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(27) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(35) XOR rng_hi_input(40) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(60) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(61) <= rng_lo_input(1) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(21) XOR rng_lo_input(26) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(35) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(42) XOR rng_lo_input(46) XOR rng_lo_input(53) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(32) XOR rng_hi_input(36) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(44) XOR rng_hi_input(46) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_lo_output(62) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(9) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(40) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(52) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(2) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(9) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(18) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(36) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(44) XOR rng_hi_input(46) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(57) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_lo_output(63) <= rng_lo_input(0) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(12) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(21) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(40) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(60) XOR rng_lo_input(62) XOR rng_hi_input(3) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(13) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(23) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(29) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(36) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(46) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(53) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(0) <= rng_lo_input(0) XOR rng_lo_input(3) XOR rng_lo_input(8) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(27) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(41) XOR rng_lo_input(43) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(4) XOR rng_hi_input(9) XOR rng_hi_input(11) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(21) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(56) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_hi_output(1) <= rng_lo_input(0) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(11) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(31) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(2) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(17) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(44) XOR rng_hi_input(48) XOR rng_hi_input(51) XOR rng_hi_input(53) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_hi_output(2) <= rng_lo_input(3) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(18) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(38) XOR rng_lo_input(41) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(25) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(43) XOR rng_hi_input(46) XOR rng_hi_input(49) XOR rng_hi_input(52) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(63);
rng_hi_output(3) <= rng_lo_input(2) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(19) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(39) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(57);
rng_hi_output(4) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(13) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(27) XOR rng_lo_input(29) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(39) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(6) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(14) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(25) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_hi_output(5) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(41) XOR rng_lo_input(47) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(54) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(42) XOR rng_hi_input(48) XOR rng_hi_input(50) XOR rng_hi_input(54) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(62);
rng_hi_output(6) <= rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(22) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(36) XOR rng_hi_input(39) XOR rng_hi_input(42) XOR rng_hi_input(48) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(58) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(7) <= rng_lo_input(0) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(22) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(63) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(11) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(55) XOR rng_hi_input(58) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(8) <= rng_lo_input(3) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(12) XOR rng_lo_input(16) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(39) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(58) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(17) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(38) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(45) XOR rng_hi_input(47) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(9) <= rng_lo_input(2) XOR rng_lo_input(5) XOR rng_lo_input(8) XOR rng_lo_input(11) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(33) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(39) XOR rng_lo_input(41) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(53) XOR rng_lo_input(56) XOR rng_lo_input(61) XOR rng_hi_input(2) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(10) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(21) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(46) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(55) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_hi_output(10) <= rng_lo_input(1) XOR rng_lo_input(3) XOR rng_lo_input(8) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(13) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(38) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(34) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(45) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(61) XOR rng_hi_input(63);
rng_hi_output(11) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(8) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(35) XOR rng_lo_input(37) XOR rng_lo_input(41) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_hi_input(0) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(30) XOR rng_hi_input(33) XOR rng_hi_input(36) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(56) XOR rng_hi_input(59) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(12) <= rng_lo_input(3) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(21) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(34) XOR rng_lo_input(40) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(51) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(61) XOR rng_hi_input(0) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(25) XOR rng_hi_input(28) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(43) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(53) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(58) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_hi_output(13) <= rng_lo_input(0) XOR rng_lo_input(3) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(50) XOR rng_lo_input(56) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_hi_input(0) XOR rng_hi_input(3) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(9) XOR rng_hi_input(13) XOR rng_hi_input(19) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(31) XOR rng_hi_input(35) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(44) XOR rng_hi_input(47) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(55) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_hi_output(14) <= rng_lo_input(1) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(29) XOR rng_lo_input(33) XOR rng_lo_input(38) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(49) XOR rng_lo_input(52) XOR rng_lo_input(56) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(10) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(41) XOR rng_hi_input(45) XOR rng_hi_input(47) XOR rng_hi_input(50) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(56) XOR rng_hi_input(59) XOR rng_hi_input(62);
rng_hi_output(15) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(10) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(22) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(27) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(37) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(47) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(56) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(60);
rng_hi_output(16) <= rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(9) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(56) XOR rng_lo_input(60) XOR rng_lo_input(63) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(5) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(12) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(46) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(55) XOR rng_hi_input(60) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(17) <= rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(17) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(27) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(40) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(7) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(37) XOR rng_hi_input(45) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(58) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(63);
rng_hi_output(18) <= rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(11) XOR rng_lo_input(14) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(29) XOR rng_lo_input(32) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(40) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(60) XOR rng_hi_input(0) XOR rng_hi_input(2) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(10) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(46) XOR rng_hi_input(48) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(60) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(19) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(58) XOR rng_hi_input(0) XOR rng_hi_input(4) XOR rng_hi_input(7) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(35) XOR rng_hi_input(38) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(49) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_hi_output(20) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(7) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(48) XOR rng_lo_input(50) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(30) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(43) XOR rng_hi_input(48) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(61);
rng_hi_output(21) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(8) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(19) XOR rng_lo_input(21) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(31) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(45) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(17) XOR rng_hi_input(21) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(38) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(44) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(53) XOR rng_hi_input(55) XOR rng_hi_input(58) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(22) <= rng_lo_input(0) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(39) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(20) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(38) XOR rng_hi_input(45) XOR rng_hi_input(48) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(56) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_hi_output(23) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(4) XOR rng_lo_input(16) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(46) XOR rng_lo_input(53) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(10) XOR rng_hi_input(13) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(21) XOR rng_hi_input(23) XOR rng_hi_input(25) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(46) XOR rng_hi_input(49) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(62);
rng_hi_output(24) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(46) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(58) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(16) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(46) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_hi_output(25) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(18) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(46) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(59) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(14) XOR rng_hi_input(17) XOR rng_hi_input(20) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(33) XOR rng_hi_input(38) XOR rng_hi_input(40) XOR rng_hi_input(44) XOR rng_hi_input(46) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(62);
rng_hi_output(26) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(4) XOR rng_hi_input(6) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(56) XOR rng_hi_input(59) XOR rng_hi_input(63);
rng_hi_output(27) <= rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(20) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(48) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(62) XOR rng_hi_input(0) XOR rng_hi_input(2) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(51) XOR rng_hi_input(53) XOR rng_hi_input(55) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(60);
rng_hi_output(28) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(57) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(25) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(39) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(52) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_hi_output(29) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(12) XOR rng_lo_input(17) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(43) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(60) XOR rng_hi_input(0) XOR rng_hi_input(2) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(30) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(60);
rng_hi_output(30) <= rng_lo_input(6) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(34) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(31) <= rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(4) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(13) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(31) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(47) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(54) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(60);
rng_hi_output(32) <= rng_lo_input(2) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(21) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(46) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(12) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(36) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(51) XOR rng_hi_input(56) XOR rng_hi_input(59) XOR rng_hi_input(60);
rng_hi_output(33) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(10) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(29) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(38) XOR rng_lo_input(41) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(7) XOR rng_hi_input(9) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(22) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(35) XOR rng_hi_input(37) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(63);
rng_hi_output(34) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(4) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(37) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(49) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(63) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(8) XOR rng_hi_input(12) XOR rng_hi_input(15) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(32) XOR rng_hi_input(35) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(55) XOR rng_hi_input(57) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(35) <= rng_lo_input(0) XOR rng_lo_input(2) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(40) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(57) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_hi_input(0) XOR rng_hi_input(2) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(27) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(58) XOR rng_hi_input(59);
rng_hi_output(36) <= rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(42) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(49) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(62) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(31) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(48) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(60) XOR rng_hi_input(63);
rng_hi_output(37) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(27) XOR rng_lo_input(29) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(41) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(19) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(31) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(47) XOR rng_hi_input(50) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(63);
rng_hi_output(38) <= rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(25) XOR rng_lo_input(27) XOR rng_lo_input(29) XOR rng_lo_input(32) XOR rng_lo_input(35) XOR rng_lo_input(38) XOR rng_lo_input(41) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(23) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(44) XOR rng_hi_input(46) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(39) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(9) XOR rng_lo_input(11) XOR rng_lo_input(13) XOR rng_lo_input(16) XOR rng_lo_input(19) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(56) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(56) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(61);
rng_hi_output(40) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(6) XOR rng_lo_input(10) XOR rng_lo_input(12) XOR rng_lo_input(15) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(39) XOR rng_lo_input(42) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(53) XOR rng_lo_input(56) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(31) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(46) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(41) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(50) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_hi_input(0) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(13) XOR rng_hi_input(16) XOR rng_hi_input(21) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_hi_output(42) <= rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(22) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(34) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(45) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(10) XOR rng_hi_input(13) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(35) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(47) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(43) <= rng_lo_input(0) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(11) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(58) XOR rng_lo_input(61) XOR rng_hi_input(0) XOR rng_hi_input(3) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(14) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(45) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(60) XOR rng_hi_input(62);
rng_hi_output(44) <= rng_lo_input(1) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(17) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(32) XOR rng_lo_input(36) XOR rng_lo_input(40) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(11) XOR rng_hi_input(16) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(47) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(55) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(62);
rng_hi_output(45) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(9) XOR rng_lo_input(11) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(53) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(59) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(10) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(61);
rng_hi_output(46) <= rng_lo_input(0) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(9) XOR rng_lo_input(11) XOR rng_lo_input(13) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(35) XOR rng_lo_input(37) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(30) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_hi_output(47) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(9) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(52) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(44) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(56) XOR rng_hi_input(58) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(48) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(8) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(36) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(50) XOR rng_lo_input(58) XOR rng_lo_input(60) XOR rng_lo_input(62) XOR rng_hi_input(0) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(10) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(42) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(60) XOR rng_hi_input(63);
rng_hi_output(49) <= rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(29) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(46) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(49) XOR rng_hi_input(53) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_hi_output(50) <= rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(29) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(34) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(49) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(58) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(15) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(46) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(60) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(51) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(20) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(37) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(14) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(32) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(58) XOR rng_hi_input(59);
rng_hi_output(52) <= rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(12) XOR rng_lo_input(18) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(43) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(57) XOR rng_lo_input(59) XOR rng_lo_input(61) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(8) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(45) XOR rng_hi_input(46) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(53) <= rng_lo_input(0) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(7) XOR rng_lo_input(9) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(17) XOR rng_lo_input(20) XOR rng_lo_input(22) XOR rng_lo_input(25) XOR rng_lo_input(30) XOR rng_lo_input(36) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(52) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(58) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(4) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(15) XOR rng_hi_input(21) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(38) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(47) XOR rng_hi_input(49) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(62);
rng_hi_output(54) <= rng_lo_input(1) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(45) XOR rng_lo_input(48) XOR rng_lo_input(52) XOR rng_lo_input(55) XOR rng_lo_input(57) XOR rng_lo_input(60) XOR rng_lo_input(63) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(11) XOR rng_hi_input(14) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(24) XOR rng_hi_input(25) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(37) XOR rng_hi_input(41) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(50) XOR rng_hi_input(52) XOR rng_hi_input(58) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(55) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(14) XOR rng_lo_input(18) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(34) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(60) XOR rng_lo_input(62) XOR rng_hi_input(0) XOR rng_hi_input(4) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(21) XOR rng_hi_input(23) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(33) XOR rng_hi_input(36) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(54) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(61);
rng_hi_output(56) <= rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(16) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(37) XOR rng_lo_input(40) XOR rng_lo_input(42) XOR rng_lo_input(45) XOR rng_lo_input(48) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(55) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_hi_input(3) XOR rng_hi_input(6) XOR rng_hi_input(8) XOR rng_hi_input(10) XOR rng_hi_input(12) XOR rng_hi_input(15) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(33) XOR rng_hi_input(36) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(47) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(57) <= rng_lo_input(0) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(10) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(14) XOR rng_lo_input(15) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(25) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(34) XOR rng_lo_input(36) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(44) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(52) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(61) XOR rng_hi_input(0) XOR rng_hi_input(2) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(61) XOR rng_hi_input(62);
rng_hi_output(58) <= rng_lo_input(0) XOR rng_lo_input(2) XOR rng_lo_input(4) XOR rng_lo_input(7) XOR rng_lo_input(11) XOR rng_lo_input(12) XOR rng_lo_input(13) XOR rng_lo_input(14) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(37) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(43) XOR rng_lo_input(44) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(52) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(1) XOR rng_hi_input(5) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(31) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(40) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(47) XOR rng_hi_input(50) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(56) XOR rng_hi_input(60);
rng_hi_output(59) <= rng_lo_input(0) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(4) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(10) XOR rng_lo_input(16) XOR rng_lo_input(19) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(23) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(39) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(45) XOR rng_lo_input(47) XOR rng_lo_input(48) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(4) XOR rng_hi_input(6) XOR rng_hi_input(9) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(13) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(19) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(22) XOR rng_hi_input(24) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(31) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(40) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(43) XOR rng_hi_input(46) XOR rng_hi_input(51) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(61) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(60) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(5) XOR rng_lo_input(6) XOR rng_lo_input(7) XOR rng_lo_input(12) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(20) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(26) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(35) XOR rng_lo_input(37) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(46) XOR rng_lo_input(49) XOR rng_lo_input(51) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_lo_input(63) XOR rng_hi_input(0) XOR rng_hi_input(2) XOR rng_hi_input(3) XOR rng_hi_input(5) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(12) XOR rng_hi_input(14) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(20) XOR rng_hi_input(24) XOR rng_hi_input(26) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(43) XOR rng_hi_input(44) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(58) XOR rng_hi_input(59);
rng_hi_output(61) <= rng_lo_input(0) XOR rng_lo_input(1) XOR rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(10) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(24) XOR rng_lo_input(27) XOR rng_lo_input(28) XOR rng_lo_input(30) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(35) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(38) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(43) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(48) XOR rng_lo_input(49) XOR rng_lo_input(50) XOR rng_lo_input(51) XOR rng_lo_input(52) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(60) XOR rng_lo_input(62) XOR rng_hi_input(0) XOR rng_hi_input(1) XOR rng_hi_input(2) XOR rng_hi_input(6) XOR rng_hi_input(7) XOR rng_hi_input(11) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(20) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(25) XOR rng_hi_input(26) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(32) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(39) XOR rng_hi_input(41) XOR rng_hi_input(42) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(48) XOR rng_hi_input(49) XOR rng_hi_input(51) XOR rng_hi_input(56) XOR rng_hi_input(57) XOR rng_hi_input(59) XOR rng_hi_input(61);
rng_hi_output(62) <= rng_lo_input(2) XOR rng_lo_input(3) XOR rng_lo_input(5) XOR rng_lo_input(7) XOR rng_lo_input(8) XOR rng_lo_input(9) XOR rng_lo_input(13) XOR rng_lo_input(16) XOR rng_lo_input(17) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(23) XOR rng_lo_input(24) XOR rng_lo_input(25) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(32) XOR rng_lo_input(36) XOR rng_lo_input(37) XOR rng_lo_input(39) XOR rng_lo_input(40) XOR rng_lo_input(41) XOR rng_lo_input(42) XOR rng_lo_input(43) XOR rng_lo_input(46) XOR rng_lo_input(51) XOR rng_lo_input(53) XOR rng_lo_input(54) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(58) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_hi_input(4) XOR rng_hi_input(6) XOR rng_hi_input(11) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(18) XOR rng_hi_input(22) XOR rng_hi_input(23) XOR rng_hi_input(25) XOR rng_hi_input(27) XOR rng_hi_input(29) XOR rng_hi_input(30) XOR rng_hi_input(33) XOR rng_hi_input(35) XOR rng_hi_input(36) XOR rng_hi_input(37) XOR rng_hi_input(41) XOR rng_hi_input(43) XOR rng_hi_input(50) XOR rng_hi_input(51) XOR rng_hi_input(52) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(62) XOR rng_hi_input(63);
rng_hi_output(63) <= rng_lo_input(0) XOR rng_lo_input(2) XOR rng_lo_input(4) XOR rng_lo_input(6) XOR rng_lo_input(8) XOR rng_lo_input(15) XOR rng_lo_input(16) XOR rng_lo_input(18) XOR rng_lo_input(20) XOR rng_lo_input(21) XOR rng_lo_input(22) XOR rng_lo_input(25) XOR rng_lo_input(28) XOR rng_lo_input(29) XOR rng_lo_input(30) XOR rng_lo_input(31) XOR rng_lo_input(32) XOR rng_lo_input(33) XOR rng_lo_input(34) XOR rng_lo_input(37) XOR rng_lo_input(40) XOR rng_lo_input(43) XOR rng_lo_input(45) XOR rng_lo_input(46) XOR rng_lo_input(52) XOR rng_lo_input(55) XOR rng_lo_input(56) XOR rng_lo_input(57) XOR rng_lo_input(59) XOR rng_lo_input(60) XOR rng_lo_input(61) XOR rng_lo_input(62) XOR rng_hi_input(1) XOR rng_hi_input(3) XOR rng_hi_input(4) XOR rng_hi_input(7) XOR rng_hi_input(8) XOR rng_hi_input(10) XOR rng_hi_input(11) XOR rng_hi_input(12) XOR rng_hi_input(15) XOR rng_hi_input(16) XOR rng_hi_input(17) XOR rng_hi_input(20) XOR rng_hi_input(21) XOR rng_hi_input(24) XOR rng_hi_input(27) XOR rng_hi_input(28) XOR rng_hi_input(29) XOR rng_hi_input(32) XOR rng_hi_input(34) XOR rng_hi_input(35) XOR rng_hi_input(37) XOR rng_hi_input(38) XOR rng_hi_input(39) XOR rng_hi_input(40) XOR rng_hi_input(42) XOR rng_hi_input(46) XOR rng_hi_input(47) XOR rng_hi_input(49) XOR rng_hi_input(50) XOR rng_hi_input(53) XOR rng_hi_input(54) XOR rng_hi_input(55) XOR rng_hi_input(57) XOR rng_hi_input(58) XOR rng_hi_input(59) XOR rng_hi_input(60) XOR rng_hi_input(61) XOR rng_hi_input(62);

END arch;